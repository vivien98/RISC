--initialize t3 with 111